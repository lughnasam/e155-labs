module lab3_lm(input logic reset,
               input logic [3:0] rows, cols,
               output logic [6:0] segout,
               output logic lpwr, rpwr);

    logic [3:0] cur_in, cur_num, prev_num;


    synchronizer (.WIDTH(4)) 

endmodule